
`ifndef APB_SVH
`define APB_SVH


`include "apb_transfer.sv"
`include "apb_config.sv"

`include "apb_master_driver.svh"
`include "apb_master_monitor.svh"
`include "apb_master_sequencer.svh"
`include "apb_master_agent.svh"

// `include "apb_slave_driver.svh"
// `include "apb_slave_monitor.svh"
// `include "apb_slave_sequencer.svh"
// `include "apb_slave_agent.svh"


`include "apb_master_driver.sv"       
`include "apb_master_monitor.sv"
`include "apb_master_sequencer.sv"
`include "apb_master_agent.sv"
`include "apb_master_seq_lib.sv"

// `include "apb_slave_driver.sv"       
// `include "apb_slave_monitor.sv"
// `include "apb_slave_sequencer.sv"
// `include "apb_slave_agent.sv"
// `include "apb_slave_seq_lib.sv"



   
`endif //  `ifndef APB_SVH
